-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 5
entity work_outputs_t_to_bytes_0CLK_82755757 is
port(
 x : in work_outputs_t;
 return_output : out uint8_t_array_4_t);
end work_outputs_t_to_bytes_0CLK_82755757;
architecture arch of work_outputs_t_to_bytes_0CLK_82755757 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes[work_outputs_t_bytes_t_h_l19_c40_821d]
signal FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x : signed(7 downto 0);
signal FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output : uint8_t_array_1_t;

-- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes[work_outputs_t_bytes_t_h_l19_c40_821d]
signal FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x : signed(7 downto 0);
signal FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output : uint8_t_array_1_t;

-- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes[work_outputs_t_bytes_t_h_l19_c40_821d]
signal FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x : signed(7 downto 0);
signal FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output : uint8_t_array_1_t;

-- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes[work_outputs_t_bytes_t_h_l19_c40_821d]
signal FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x : signed(7 downto 0);
signal FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output : uint8_t_array_1_t;

function CONST_REF_RD_uint8_t_array_4_t_uint8_t_array_4_t_4a68( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned) return uint8_t_array_4_t is
 
  variable base : uint8_t_array_4_t; 
  variable return_output : uint8_t_array_4_t;
begin
      base.data(0) := ref_toks_0;
      base.data(1) := ref_toks_1;
      base.data(2) := ref_toks_2;
      base.data(3) := ref_toks_3;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d : 0 clocks latency
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d : entity work.int8_t_to_bytes_0CLK_23f04728 port map (
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x,
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output);

-- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d : 0 clocks latency
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d : entity work.int8_t_to_bytes_0CLK_23f04728 port map (
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x,
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output);

-- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d : 0 clocks latency
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d : entity work.int8_t_to_bytes_0CLK_23f04728 port map (
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x,
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output);

-- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d : 0 clocks latency
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d : entity work.int8_t_to_bytes_0CLK_23f04728 port map (
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x,
FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 x,
 -- All submodule outputs
 FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output,
 FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output,
 FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output,
 FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : uint8_t_array_4_t;
 variable VAR_x : work_outputs_t;
 variable VAR_rv : uint8_t_array_4_t;
 variable VAR_pos : unsigned(2 downto 0);
 variable VAR_field_pos : unsigned(2 downto 0);
 variable VAR_result_dim_0 : unsigned(1 downto 0);
 variable VAR_result_dim_1 : unsigned(1 downto 0);
 variable VAR_result_elem_bytes : uint8_t_array_1_t;
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x : signed(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_CONST_REF_RD_int8_t_work_outputs_t_result_0_0_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output : signed(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x : signed(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_CONST_REF_RD_int8_t_work_outputs_t_result_0_1_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output : signed(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x : signed(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_CONST_REF_RD_int8_t_work_outputs_t_result_1_0_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output : signed(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x : signed(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_CONST_REF_RD_int8_t_work_outputs_t_result_1_1_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output : signed(7 downto 0);
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_4_t_uint8_t_array_4_t_4a68_work_outputs_t_bytes_t_h_l28_c12_f253_return_output : uint8_t_array_4_t;
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_x := x;

     -- Submodule level 0
     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_CONST_REF_RD_int8_t_work_outputs_t_result_0_1_d41d[work_outputs_t_bytes_t_h_l19_c56_763f] LATENCY=0
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_CONST_REF_RD_int8_t_work_outputs_t_result_0_1_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output := VAR_x.result(0)(1);

     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_CONST_REF_RD_int8_t_work_outputs_t_result_1_0_d41d[work_outputs_t_bytes_t_h_l19_c56_763f] LATENCY=0
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_CONST_REF_RD_int8_t_work_outputs_t_result_1_0_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output := VAR_x.result(1)(0);

     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_CONST_REF_RD_int8_t_work_outputs_t_result_0_0_d41d[work_outputs_t_bytes_t_h_l19_c56_763f] LATENCY=0
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_CONST_REF_RD_int8_t_work_outputs_t_result_0_0_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output := VAR_x.result(0)(0);

     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_CONST_REF_RD_int8_t_work_outputs_t_result_1_1_d41d[work_outputs_t_bytes_t_h_l19_c56_763f] LATENCY=0
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_CONST_REF_RD_int8_t_work_outputs_t_result_1_1_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output := VAR_x.result(1)(1);

     -- Submodule level 1
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x := VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_CONST_REF_RD_int8_t_work_outputs_t_result_0_0_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output;
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x := VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_CONST_REF_RD_int8_t_work_outputs_t_result_0_1_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output;
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x := VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_CONST_REF_RD_int8_t_work_outputs_t_result_1_0_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output;
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x := VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_CONST_REF_RD_int8_t_work_outputs_t_result_1_1_d41d_work_outputs_t_bytes_t_h_l19_c56_763f_return_output;
     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes[work_outputs_t_bytes_t_h_l19_c40_821d] LATENCY=0
     -- Inputs
     FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x <= VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x;
     -- Outputs
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output := FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output;

     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes[work_outputs_t_bytes_t_h_l19_c40_821d] LATENCY=0
     -- Inputs
     FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x <= VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x;
     -- Outputs
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output := FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output;

     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes[work_outputs_t_bytes_t_h_l19_c40_821d] LATENCY=0
     -- Inputs
     FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x <= VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x;
     -- Outputs
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output := FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output;

     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes[work_outputs_t_bytes_t_h_l19_c40_821d] LATENCY=0
     -- Inputs
     FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x <= VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_x;
     -- Outputs
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output := FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output;

     -- Submodule level 2
     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d[work_outputs_t_bytes_t_h_l22_c20_011c] LATENCY=0
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output := VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output.data(0);

     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d[work_outputs_t_bytes_t_h_l22_c20_011c] LATENCY=0
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output := VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output.data(0);

     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d[work_outputs_t_bytes_t_h_l22_c20_011c] LATENCY=0
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output := VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output.data(0);

     -- FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d[work_outputs_t_bytes_t_h_l22_c20_011c] LATENCY=0
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output := VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_int8_t_to_bytes_work_outputs_t_bytes_t_h_l19_c40_821d_return_output.data(0);

     -- Submodule level 3
     -- CONST_REF_RD_uint8_t_array_4_t_uint8_t_array_4_t_4a68[work_outputs_t_bytes_t_h_l28_c12_f253] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_4_t_uint8_t_array_4_t_4a68_work_outputs_t_bytes_t_h_l28_c12_f253_return_output := CONST_REF_RD_uint8_t_array_4_t_uint8_t_array_4_t_4a68(
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output,
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_0_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output,
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_0_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output,
     VAR_FOR_work_outputs_t_bytes_t_h_l16_c1_c8e1_ITER_1_FOR_work_outputs_t_bytes_t_h_l18_c1_7320_ITER_1_FOR_work_outputs_t_bytes_t_h_l20_c2_3c02_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_1_t_data_0_d41d_work_outputs_t_bytes_t_h_l22_c20_011c_return_output);

     -- Submodule level 4
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_4_t_uint8_t_array_4_t_4a68_work_outputs_t_bytes_t_h_l28_c12_f253_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
