-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 19
entity skid_buf_rmii_eth_mac_tx_fifo_0CLK_83e31706 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 stream_in : in axis8_t_stream_t;
 ready_for_stream_out : in unsigned(0 downto 0);
 return_output : out skid_buf_rmii_eth_mac_tx_fifo_t);
end skid_buf_rmii_eth_mac_tx_fifo_0CLK_83e31706;
architecture arch of skid_buf_rmii_eth_mac_tx_fifo_0CLK_83e31706 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal buff : axis8_t_stream_t := axis8_t_stream_t_NULL;
signal skid_buff : axis8_t_stream_t := axis8_t_stream_t_NULL;
signal output_is_skid_buff : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_buff : axis8_t_stream_t;
signal REG_COMB_skid_buff : axis8_t_stream_t;
signal REG_COMB_output_is_skid_buff : unsigned(0 downto 0);

-- Resolved maybe from input reg clock enable
signal clk_en_internal : std_logic;
-- Each function instance gets signals
-- o_MUX[rmii_eth_mac_c_l14_c681_5240]
signal o_MUX_rmii_eth_mac_c_l14_c681_5240_cond : unsigned(0 downto 0);
signal o_MUX_rmii_eth_mac_c_l14_c681_5240_iftrue : skid_buf_rmii_eth_mac_tx_fifo_t;
signal o_MUX_rmii_eth_mac_c_l14_c681_5240_iffalse : skid_buf_rmii_eth_mac_tx_fifo_t;
signal o_MUX_rmii_eth_mac_c_l14_c681_5240_return_output : skid_buf_rmii_eth_mac_tx_fifo_t;

-- UNARY_OP_NOT[rmii_eth_mac_c_l14_c757_c5fd]
signal UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_return_output : unsigned(0 downto 0);

-- UNARY_OP_NOT[rmii_eth_mac_c_l14_c822_2899]
signal UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_return_output : unsigned(0 downto 0);

-- skid_buff_MUX[rmii_eth_mac_c_l14_c841_19a1]
signal skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond : unsigned(0 downto 0);
signal skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue : axis8_t_stream_t;
signal skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse : axis8_t_stream_t;
signal skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output : axis8_t_stream_t;

-- buff_MUX[rmii_eth_mac_c_l14_c841_19a1]
signal buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond : unsigned(0 downto 0);
signal buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue : axis8_t_stream_t;
signal buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse : axis8_t_stream_t;
signal buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output : axis8_t_stream_t;

-- skid_buff_MUX[rmii_eth_mac_c_l14_c868_7779]
signal skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond : unsigned(0 downto 0);
signal skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue : axis8_t_stream_t;
signal skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse : axis8_t_stream_t;
signal skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output : axis8_t_stream_t;

-- buff_MUX[rmii_eth_mac_c_l14_c868_7779]
signal buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond : unsigned(0 downto 0);
signal buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue : axis8_t_stream_t;
signal buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse : axis8_t_stream_t;
signal buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output : axis8_t_stream_t;

-- UNARY_OP_NOT[rmii_eth_mac_c_l14_c949_bb5e]
signal UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_return_output : unsigned(0 downto 0);

-- BIN_OP_OR[rmii_eth_mac_c_l14_c949_a869]
signal BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_left : unsigned(0 downto 0);
signal BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_right : unsigned(0 downto 0);
signal BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_return_output : unsigned(0 downto 0);

-- output_is_skid_buff_MUX[rmii_eth_mac_c_l14_c945_13fb]
signal output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_cond : unsigned(0 downto 0);
signal output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue : unsigned(0 downto 0);
signal output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse : unsigned(0 downto 0);
signal output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output : unsigned(0 downto 0);

-- skid_buff_valid_MUX[rmii_eth_mac_c_l14_c945_13fb]
signal skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond : unsigned(0 downto 0);
signal skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue : unsigned(0 downto 0);
signal skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse : unsigned(0 downto 0);
signal skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output : unsigned(0 downto 0);

-- buff_valid_MUX[rmii_eth_mac_c_l14_c945_13fb]
signal buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond : unsigned(0 downto 0);
signal buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue : unsigned(0 downto 0);
signal buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse : unsigned(0 downto 0);
signal buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output : unsigned(0 downto 0);

-- skid_buff_valid_MUX[rmii_eth_mac_c_l14_c993_c374]
signal skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond : unsigned(0 downto 0);
signal skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue : unsigned(0 downto 0);
signal skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse : unsigned(0 downto 0);
signal skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output : unsigned(0 downto 0);

-- buff_valid_MUX[rmii_eth_mac_c_l14_c993_c374]
signal buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond : unsigned(0 downto 0);
signal buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue : unsigned(0 downto 0);
signal buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse : unsigned(0 downto 0);
signal buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output : unsigned(0 downto 0);

-- UNARY_OP_NOT[rmii_eth_mac_c_l14_c1087_be7c]
signal UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_return_output : unsigned(0 downto 0);

function CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3( ref_toks_0 : axis8_t_stream_t;
 ref_toks_1 : unsigned) return skid_buf_rmii_eth_mac_tx_fifo_t is
 
  variable base : skid_buf_rmii_eth_mac_tx_fifo_t; 
  variable return_output : skid_buf_rmii_eth_mac_tx_fifo_t;
begin
      base.stream_out := ref_toks_0;
      base.ready_for_stream_in := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee( ref_toks_0 : axis8_t_stream_t;
 ref_toks_1 : unsigned) return axis8_t_stream_t is
 
  variable base : axis8_t_stream_t; 
  variable return_output : axis8_t_stream_t;
begin
      base := ref_toks_0;
      base.valid := ref_toks_1;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- o_MUX_rmii_eth_mac_c_l14_c681_5240 : 0 clocks latency
o_MUX_rmii_eth_mac_c_l14_c681_5240 : entity work.MUX_uint1_t_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_0CLK_de264c78 port map (
o_MUX_rmii_eth_mac_c_l14_c681_5240_cond,
o_MUX_rmii_eth_mac_c_l14_c681_5240_iftrue,
o_MUX_rmii_eth_mac_c_l14_c681_5240_iffalse,
o_MUX_rmii_eth_mac_c_l14_c681_5240_return_output);

-- UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd : 0 clocks latency
UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_expr,
UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_return_output);

-- UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899 : 0 clocks latency
UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_expr,
UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_return_output);

-- skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1 : 0 clocks latency
skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1 : entity work.MUX_uint1_t_axis8_t_stream_t_axis8_t_stream_t_0CLK_de264c78 port map (
skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond,
skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue,
skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse,
skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output);

-- buff_MUX_rmii_eth_mac_c_l14_c841_19a1 : 0 clocks latency
buff_MUX_rmii_eth_mac_c_l14_c841_19a1 : entity work.MUX_uint1_t_axis8_t_stream_t_axis8_t_stream_t_0CLK_de264c78 port map (
buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond,
buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue,
buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse,
buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output);

-- skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779 : 0 clocks latency
skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779 : entity work.MUX_uint1_t_axis8_t_stream_t_axis8_t_stream_t_0CLK_de264c78 port map (
skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond,
skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue,
skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse,
skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output);

-- buff_MUX_rmii_eth_mac_c_l14_c868_7779 : 0 clocks latency
buff_MUX_rmii_eth_mac_c_l14_c868_7779 : entity work.MUX_uint1_t_axis8_t_stream_t_axis8_t_stream_t_0CLK_de264c78 port map (
buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond,
buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue,
buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse,
buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output);

-- UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e : 0 clocks latency
UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_expr,
UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_return_output);

-- BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869 : 0 clocks latency
BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869 : entity work.BIN_OP_OR_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_left,
BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_right,
BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_return_output);

-- output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb : 0 clocks latency
output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_cond,
output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue,
output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse,
output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output);

-- skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb : 0 clocks latency
skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond,
skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue,
skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse,
skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output);

-- buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb : 0 clocks latency
buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond,
buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue,
buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse,
buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output);

-- skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374 : 0 clocks latency
skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond,
skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue,
skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse,
skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output);

-- buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374 : 0 clocks latency
buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond,
buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue,
buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse,
buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output);

-- UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c : 0 clocks latency
UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_expr,
UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_return_output);



-- Resolve what clock enable to use for user logic
clk_en_internal <= CLOCK_ENABLE(0);
-- Combinatorial process for pipeline stages
process (
CLOCK_ENABLE,
clk_en_internal,
 -- Inputs
 stream_in,
 ready_for_stream_out,
 -- Registers
 buff,
 skid_buff,
 output_is_skid_buff,
 -- All submodule outputs
 o_MUX_rmii_eth_mac_c_l14_c681_5240_return_output,
 UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_return_output,
 UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_return_output,
 skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output,
 buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output,
 skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output,
 buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output,
 UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_return_output,
 BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_return_output,
 output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output,
 skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output,
 buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output,
 skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output,
 buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output,
 UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : skid_buf_rmii_eth_mac_tx_fifo_t;
 variable VAR_stream_in : axis8_t_stream_t;
 variable VAR_ready_for_stream_out : unsigned(0 downto 0);
 variable VAR_o : skid_buf_rmii_eth_mac_tx_fifo_t;
 variable VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_iftrue : skid_buf_rmii_eth_mac_tx_fifo_t;
 variable VAR_o_TRUE_INPUT_MUX_CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3_rmii_eth_mac_c_l14_c681_5240_return_output : skid_buf_rmii_eth_mac_tx_fifo_t;
 variable VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_iffalse : skid_buf_rmii_eth_mac_tx_fifo_t;
 variable VAR_o_FALSE_INPUT_MUX_CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3_rmii_eth_mac_c_l14_c681_5240_return_output : skid_buf_rmii_eth_mac_tx_fifo_t;
 variable VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_return_output : skid_buf_rmii_eth_mac_tx_fifo_t;
 variable VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_c757_a861_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_c822_a9cf_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_skid_buf_rmii_eth_mac_tx_fifo_t_ready_for_stream_in_d41d_rmii_eth_mac_c_l14_c844_d31a_return_output : unsigned(0 downto 0);
 variable VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue : axis8_t_stream_t;
 variable VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output : axis8_t_stream_t;
 variable VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse : axis8_t_stream_t;
 variable VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output : axis8_t_stream_t;
 variable VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond : unsigned(0 downto 0);
 variable VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue : axis8_t_stream_t;
 variable VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output : axis8_t_stream_t;
 variable VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse : axis8_t_stream_t;
 variable VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output : axis8_t_stream_t;
 variable VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond : unsigned(0 downto 0);
 variable VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue : axis8_t_stream_t;
 variable VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse : axis8_t_stream_t;
 variable VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond : unsigned(0 downto 0);
 variable VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue : axis8_t_stream_t;
 variable VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse : axis8_t_stream_t;
 variable VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_skid_buf_rmii_eth_mac_tx_fifo_t_stream_out_valid_d41d_rmii_eth_mac_c_l14_c949_53c2_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_return_output : unsigned(0 downto 0);
 variable VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue : unsigned(0 downto 0);
 variable VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse : unsigned(0 downto 0);
 variable VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output : unsigned(0 downto 0);
 variable VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_cond : unsigned(0 downto 0);
 variable VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue : unsigned(0 downto 0);
 variable VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output : unsigned(0 downto 0);
 variable VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse : unsigned(0 downto 0);
 variable VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output : unsigned(0 downto 0);
 variable VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond : unsigned(0 downto 0);
 variable VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue : unsigned(0 downto 0);
 variable VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output : unsigned(0 downto 0);
 variable VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse : unsigned(0 downto 0);
 variable VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output : unsigned(0 downto 0);
 variable VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond : unsigned(0 downto 0);
 variable VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue : unsigned(0 downto 0);
 variable VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse : unsigned(0 downto 0);
 variable VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond : unsigned(0 downto 0);
 variable VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue : unsigned(0 downto 0);
 variable VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse : unsigned(0 downto 0);
 variable VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_return_output : unsigned(0 downto 0);
 variable VAR_buff_CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee_rmii_eth_mac_c_l14_c455_0664_return_output : axis8_t_stream_t;
 variable VAR_skid_buff_CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee_rmii_eth_mac_c_l14_c455_0664_return_output : axis8_t_stream_t;
 variable VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_DUPLICATE_7662_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_DUPLICATE_8c0f_return_output : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_buff : axis8_t_stream_t;
variable REG_VAR_skid_buff : axis8_t_stream_t;
variable REG_VAR_output_is_skid_buff : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_buff := buff;
  REG_VAR_skid_buff := skid_buff;
  REG_VAR_output_is_skid_buff := output_is_skid_buff;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue := to_unsigned(0, 1);
     VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE(0) := clk_en_internal;
     -- Mux in inputs
     VAR_stream_in := stream_in;
     VAR_ready_for_stream_out := ready_for_stream_out;

     -- Submodule level 0
     VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse := buff;
     VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse := buff;
     VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_expr := output_is_skid_buff;
     VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond := output_is_skid_buff;
     VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond := output_is_skid_buff;
     VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_cond := output_is_skid_buff;
     VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse := output_is_skid_buff;
     VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond := output_is_skid_buff;
     VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond := output_is_skid_buff;
     VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_right := VAR_ready_for_stream_out;
     VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse := skid_buff;
     VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue := skid_buff;
     VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue := VAR_stream_in;
     VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse := VAR_stream_in;
     -- skid_buff_MUX[rmii_eth_mac_c_l14_c868_7779] LATENCY=0
     -- Inputs
     skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond <= VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond;
     skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue <= VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue;
     skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse <= VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse;
     -- Outputs
     VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output := skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output;

     -- buff_MUX[rmii_eth_mac_c_l14_c868_7779] LATENCY=0
     -- Inputs
     buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond <= VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_cond;
     buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue <= VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iftrue;
     buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse <= VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_iffalse;
     -- Outputs
     VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output := buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output;

     -- CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d[rmii_eth_mac_c_l14_c757_a861] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_c757_a861_return_output := buff.valid;

     -- CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d[rmii_eth_mac_c_l14_c822_a9cf] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_c822_a9cf_return_output := skid_buff.valid;

     -- UNARY_OP_NOT[rmii_eth_mac_c_l14_c1087_be7c] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_expr <= VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_return_output := UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_return_output;

     -- Submodule level 1
     VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_expr := VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_c757_a861_return_output;
     VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_expr := VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_c822_a9cf_return_output;
     VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue := VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c1087_be7c_return_output;
     VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue := VAR_buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output;
     VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue := VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c868_7779_return_output;
     -- UNARY_OP_NOT[rmii_eth_mac_c_l14_c757_c5fd] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_expr <= VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_return_output := UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_return_output;

     -- UNARY_OP_NOT[rmii_eth_mac_c_l14_c822_2899] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_expr <= VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_return_output := UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_return_output;

     -- Submodule level 2
     -- o_FALSE_INPUT_MUX_CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3[rmii_eth_mac_c_l14_c681_5240] LATENCY=0
     VAR_o_FALSE_INPUT_MUX_CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3_rmii_eth_mac_c_l14_c681_5240_return_output := CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3(
     buff,
     VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c822_2899_return_output);

     -- o_TRUE_INPUT_MUX_CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3[rmii_eth_mac_c_l14_c681_5240] LATENCY=0
     VAR_o_TRUE_INPUT_MUX_CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3_rmii_eth_mac_c_l14_c681_5240_return_output := CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3(
     skid_buff,
     VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c757_c5fd_return_output);

     -- Submodule level 3
     VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_iffalse := VAR_o_FALSE_INPUT_MUX_CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3_rmii_eth_mac_c_l14_c681_5240_return_output;
     VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_iftrue := VAR_o_TRUE_INPUT_MUX_CONST_REF_RD_skid_buf_rmii_eth_mac_tx_fifo_t_skid_buf_rmii_eth_mac_tx_fifo_t_69f3_rmii_eth_mac_c_l14_c681_5240_return_output;
     -- o_MUX[rmii_eth_mac_c_l14_c681_5240] LATENCY=0
     -- Inputs
     o_MUX_rmii_eth_mac_c_l14_c681_5240_cond <= VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_cond;
     o_MUX_rmii_eth_mac_c_l14_c681_5240_iftrue <= VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_iftrue;
     o_MUX_rmii_eth_mac_c_l14_c681_5240_iffalse <= VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_iffalse;
     -- Outputs
     VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_return_output := o_MUX_rmii_eth_mac_c_l14_c681_5240_return_output;

     -- Submodule level 4
     VAR_return_output := VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_return_output;
     -- CONST_REF_RD_uint1_t_skid_buf_rmii_eth_mac_tx_fifo_t_stream_out_valid_d41d[rmii_eth_mac_c_l14_c949_53c2] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_skid_buf_rmii_eth_mac_tx_fifo_t_stream_out_valid_d41d_rmii_eth_mac_c_l14_c949_53c2_return_output := VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_return_output.stream_out.valid;

     -- CONST_REF_RD_uint1_t_skid_buf_rmii_eth_mac_tx_fifo_t_ready_for_stream_in_d41d[rmii_eth_mac_c_l14_c844_d31a] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_skid_buf_rmii_eth_mac_tx_fifo_t_ready_for_stream_in_d41d_rmii_eth_mac_c_l14_c844_d31a_return_output := VAR_o_MUX_rmii_eth_mac_c_l14_c681_5240_return_output.ready_for_stream_in;

     -- Submodule level 5
     VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond := VAR_CONST_REF_RD_uint1_t_skid_buf_rmii_eth_mac_tx_fifo_t_ready_for_stream_in_d41d_rmii_eth_mac_c_l14_c844_d31a_return_output;
     VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond := VAR_CONST_REF_RD_uint1_t_skid_buf_rmii_eth_mac_tx_fifo_t_ready_for_stream_in_d41d_rmii_eth_mac_c_l14_c844_d31a_return_output;
     VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_expr := VAR_CONST_REF_RD_uint1_t_skid_buf_rmii_eth_mac_tx_fifo_t_stream_out_valid_d41d_rmii_eth_mac_c_l14_c949_53c2_return_output;
     -- buff_MUX[rmii_eth_mac_c_l14_c841_19a1] LATENCY=0
     -- Inputs
     buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond <= VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond;
     buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue <= VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue;
     buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse <= VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse;
     -- Outputs
     VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output := buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output;

     -- skid_buff_MUX[rmii_eth_mac_c_l14_c841_19a1] LATENCY=0
     -- Inputs
     skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond <= VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_cond;
     skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue <= VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iftrue;
     skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse <= VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_iffalse;
     -- Outputs
     VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output := skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output;

     -- UNARY_OP_NOT[rmii_eth_mac_c_l14_c949_bb5e] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_expr <= VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_return_output := UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_return_output;

     -- Submodule level 6
     VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_left := VAR_UNARY_OP_NOT_rmii_eth_mac_c_l14_c949_bb5e_return_output;
     -- CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_DUPLICATE_8c0f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_DUPLICATE_8c0f_return_output := VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output.valid;

     -- CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_DUPLICATE_7662 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_DUPLICATE_7662_return_output := VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output.valid;

     -- BIN_OP_OR[rmii_eth_mac_c_l14_c949_a869] LATENCY=0
     -- Inputs
     BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_left <= VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_left;
     BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_right <= VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_right;
     -- Outputs
     VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_return_output := BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_return_output;

     -- Submodule level 7
     VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond := VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_return_output;
     VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_cond := VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_return_output;
     VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond := VAR_BIN_OP_OR_rmii_eth_mac_c_l14_c949_a869_return_output;
     VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse := VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_DUPLICATE_7662_return_output;
     VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue := VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_DUPLICATE_7662_return_output;
     VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse := VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_DUPLICATE_8c0f_return_output;
     VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse := VAR_CONST_REF_RD_uint1_t_axis8_t_stream_t_valid_d41d_rmii_eth_mac_c_l14_DUPLICATE_8c0f_return_output;
     -- skid_buff_valid_MUX[rmii_eth_mac_c_l14_c993_c374] LATENCY=0
     -- Inputs
     skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond <= VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond;
     skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue <= VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue;
     skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse <= VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse;
     -- Outputs
     VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output := skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output;

     -- buff_valid_MUX[rmii_eth_mac_c_l14_c993_c374] LATENCY=0
     -- Inputs
     buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond <= VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_cond;
     buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue <= VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iftrue;
     buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse <= VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_iffalse;
     -- Outputs
     VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output := buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output;

     -- output_is_skid_buff_MUX[rmii_eth_mac_c_l14_c945_13fb] LATENCY=0
     -- Inputs
     output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_cond <= VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_cond;
     output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue <= VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue;
     output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse <= VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse;
     -- Outputs
     VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output := output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output;

     -- Submodule level 8
     VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue := VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output;
     REG_VAR_output_is_skid_buff := VAR_output_is_skid_buff_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output;
     VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue := VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c993_c374_return_output;
     -- skid_buff_valid_MUX[rmii_eth_mac_c_l14_c945_13fb] LATENCY=0
     -- Inputs
     skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond <= VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond;
     skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue <= VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue;
     skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse <= VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse;
     -- Outputs
     VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output := skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output;

     -- buff_valid_MUX[rmii_eth_mac_c_l14_c945_13fb] LATENCY=0
     -- Inputs
     buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond <= VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_cond;
     buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue <= VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iftrue;
     buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse <= VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_iffalse;
     -- Outputs
     VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output := buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output;

     -- Submodule level 9
     -- buff_CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee[rmii_eth_mac_c_l14_c455_0664] LATENCY=0
     VAR_buff_CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee_rmii_eth_mac_c_l14_c455_0664_return_output := CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee(
     VAR_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output,
     VAR_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output);

     -- skid_buff_CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee[rmii_eth_mac_c_l14_c455_0664] LATENCY=0
     VAR_skid_buff_CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee_rmii_eth_mac_c_l14_c455_0664_return_output := CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee(
     VAR_skid_buff_MUX_rmii_eth_mac_c_l14_c841_19a1_return_output,
     VAR_skid_buff_valid_MUX_rmii_eth_mac_c_l14_c945_13fb_return_output);

     -- Submodule level 10
     REG_VAR_buff := VAR_buff_CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee_rmii_eth_mac_c_l14_c455_0664_return_output;
     REG_VAR_skid_buff := VAR_skid_buff_CONST_REF_RD_axis8_t_stream_t_axis8_t_stream_t_2dee_rmii_eth_mac_c_l14_c455_0664_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_buff <= REG_VAR_buff;
REG_COMB_skid_buff <= REG_VAR_skid_buff;
REG_COMB_output_is_skid_buff <= REG_VAR_output_is_skid_buff;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if clk_en_internal='1' then
     buff <= REG_COMB_buff;
     skid_buff <= REG_COMB_skid_buff;
     output_is_skid_buff <= REG_COMB_output_is_skid_buff;
 end if;
 end if;
end process;

end arch;
