-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 17
entity bytes_to_work_inputs_t_0CLK_5670a028 is
port(
 bytes : in uint8_t_8;
 return_output : out work_inputs_t);
end bytes_to_work_inputs_t_0CLK_5670a028;
architecture arch of bytes_to_work_inputs_t_0CLK_5670a028 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t[work_inputs_t_bytes_t_h_l69_c45_ff13]
signal FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes : uint8_t_1;
signal FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output : signed(7 downto 0);

-- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t[work_inputs_t_bytes_t_h_l69_c45_ff13]
signal FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes : uint8_t_1;
signal FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output : signed(7 downto 0);

-- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t[work_inputs_t_bytes_t_h_l69_c45_ff13]
signal FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes : uint8_t_1;
signal FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output : signed(7 downto 0);

-- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t[work_inputs_t_bytes_t_h_l69_c45_ff13]
signal FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes : uint8_t_1;
signal FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output : signed(7 downto 0);

-- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t[work_inputs_t_bytes_t_h_l83_c45_bb36]
signal FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes : uint8_t_1;
signal FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output : signed(7 downto 0);

-- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t[work_inputs_t_bytes_t_h_l83_c45_bb36]
signal FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes : uint8_t_1;
signal FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output : signed(7 downto 0);

-- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t[work_inputs_t_bytes_t_h_l83_c45_bb36]
signal FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes : uint8_t_1;
signal FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output : signed(7 downto 0);

-- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t[work_inputs_t_bytes_t_h_l83_c45_bb36]
signal FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes : uint8_t_1;
signal FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output : signed(7 downto 0);

function CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41( ref_toks_0 : unsigned) return uint8_t_array_1_t is
 
  variable base : uint8_t_array_1_t; 
  variable return_output : uint8_t_array_1_t;
begin
      base.data(0) := ref_toks_0;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_work_inputs_t_work_inputs_t_1fa3( ref_toks_0 : signed;
 ref_toks_1 : signed;
 ref_toks_2 : signed;
 ref_toks_3 : signed;
 ref_toks_4 : signed;
 ref_toks_5 : signed;
 ref_toks_6 : signed;
 ref_toks_7 : signed) return work_inputs_t is
 
  variable base : work_inputs_t; 
  variable return_output : work_inputs_t;
begin
      base.matrix0(0)(0) := ref_toks_0;
      base.matrix0(0)(1) := ref_toks_1;
      base.matrix0(1)(0) := ref_toks_2;
      base.matrix0(1)(1) := ref_toks_3;
      base.matrix1(0)(0) := ref_toks_4;
      base.matrix1(0)(1) := ref_toks_5;
      base.matrix1(1)(0) := ref_toks_6;
      base.matrix1(1)(1) := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13 : 0 clocks latency
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13 : entity work.bytes_to_int8_t_0CLK_23f04728 port map (
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes,
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output);

-- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13 : 0 clocks latency
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13 : entity work.bytes_to_int8_t_0CLK_23f04728 port map (
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes,
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output);

-- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13 : 0 clocks latency
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13 : entity work.bytes_to_int8_t_0CLK_23f04728 port map (
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes,
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output);

-- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13 : 0 clocks latency
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13 : entity work.bytes_to_int8_t_0CLK_23f04728 port map (
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes,
FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output);

-- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36 : 0 clocks latency
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36 : entity work.bytes_to_int8_t_0CLK_23f04728 port map (
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes,
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output);

-- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36 : 0 clocks latency
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36 : entity work.bytes_to_int8_t_0CLK_23f04728 port map (
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes,
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output);

-- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36 : 0 clocks latency
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36 : entity work.bytes_to_int8_t_0CLK_23f04728 port map (
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes,
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output);

-- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36 : 0 clocks latency
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36 : entity work.bytes_to_int8_t_0CLK_23f04728 port map (
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes,
FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 bytes,
 -- All submodule outputs
 FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output,
 FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output,
 FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output,
 FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output,
 FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output,
 FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output,
 FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output,
 FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : work_inputs_t;
 variable VAR_bytes : uint8_t_8;
 variable VAR_rv : work_inputs_t;
 variable VAR_pos : unsigned(3 downto 0);
 variable VAR_field_pos : unsigned(3 downto 0);
 variable VAR_matrix0_dim_0 : unsigned(1 downto 0);
 variable VAR_matrix0_dim_1 : unsigned(1 downto 0);
 variable VAR_matrix0_elem_bytes : uint8_t_array_1_t;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes : uint8_t_1;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output : signed(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes : uint8_t_1;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output : signed(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes : uint8_t_1;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output : signed(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes : uint8_t_1;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output : signed(7 downto 0);
 variable VAR_matrix1_dim_0 : unsigned(1 downto 0);
 variable VAR_matrix1_dim_1 : unsigned(1 downto 0);
 variable VAR_matrix1_elem_bytes : uint8_t_array_1_t;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes : uint8_t_1;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output : signed(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes : uint8_t_1;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output : signed(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes : uint8_t_1;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output : signed(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output : unsigned(7 downto 0);
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes : uint8_t_1;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output : uint8_t_array_1_t;
 variable VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_work_inputs_t_work_inputs_t_1fa3_work_inputs_t_bytes_t_h_l87_c12_d3f7_return_output : work_inputs_t;
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_bytes := bytes;

     -- Submodule level 0
     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d[work_inputs_t_bytes_t_h_l80_c42_a3a0] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output := VAR_bytes(6);

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d[work_inputs_t_bytes_t_h_l80_c42_a3a0] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output := VAR_bytes(7);

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d[work_inputs_t_bytes_t_h_l80_c42_a3a0] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output := VAR_bytes(4);

     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d[work_inputs_t_bytes_t_h_l66_c42_4a95] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output := VAR_bytes(3);

     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d[work_inputs_t_bytes_t_h_l66_c42_4a95] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output := VAR_bytes(1);

     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d[work_inputs_t_bytes_t_h_l66_c42_4a95] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output := VAR_bytes(2);

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d[work_inputs_t_bytes_t_h_l80_c42_a3a0] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output := VAR_bytes(5);

     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d[work_inputs_t_bytes_t_h_l66_c42_4a95] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output := VAR_bytes(0);

     -- Submodule level 1
     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41[work_inputs_t_bytes_t_h_l69_c61_4e04] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output := CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41(
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output);

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41[work_inputs_t_bytes_t_h_l83_c61_d47c] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output := CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41(
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output);

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41[work_inputs_t_bytes_t_h_l83_c61_d47c] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output := CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41(
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output);

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41[work_inputs_t_bytes_t_h_l83_c61_d47c] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output := CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41(
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output);

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41[work_inputs_t_bytes_t_h_l83_c61_d47c] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output := CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41(
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_FOR_work_inputs_t_bytes_t_h_l78_c2_f280_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_work_inputs_t_bytes_t_h_l80_c42_a3a0_return_output);

     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41[work_inputs_t_bytes_t_h_l69_c61_4e04] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output := CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41(
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output);

     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41[work_inputs_t_bytes_t_h_l69_c61_4e04] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output := CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41(
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output);

     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41[work_inputs_t_bytes_t_h_l69_c61_4e04] LATENCY=0
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output := CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41(
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_FOR_work_inputs_t_bytes_t_h_l64_c2_76ef_ITER_0_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_work_inputs_t_bytes_t_h_l66_c42_4a95_return_output);

     -- Submodule level 2
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes := VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output.data;
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes := VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output.data;
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes := VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output.data;
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes := VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l69_c61_4e04_return_output.data;
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes := VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output.data;
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes := VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output.data;
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes := VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output.data;
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes := VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_CONST_REF_RD_uint8_t_array_1_t_uint8_t_array_1_t_5b41_work_inputs_t_bytes_t_h_l83_c61_d47c_return_output.data;
     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t[work_inputs_t_bytes_t_h_l69_c45_ff13] LATENCY=0
     -- Inputs
     FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes <= VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes;
     -- Outputs
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output := FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output;

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t[work_inputs_t_bytes_t_h_l83_c45_bb36] LATENCY=0
     -- Inputs
     FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes <= VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes;
     -- Outputs
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output := FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output;

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t[work_inputs_t_bytes_t_h_l83_c45_bb36] LATENCY=0
     -- Inputs
     FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes <= VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes;
     -- Outputs
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output := FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output;

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t[work_inputs_t_bytes_t_h_l83_c45_bb36] LATENCY=0
     -- Inputs
     FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes <= VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes;
     -- Outputs
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output := FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output;

     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t[work_inputs_t_bytes_t_h_l69_c45_ff13] LATENCY=0
     -- Inputs
     FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes <= VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes;
     -- Outputs
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output := FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output;

     -- FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t[work_inputs_t_bytes_t_h_l83_c45_bb36] LATENCY=0
     -- Inputs
     FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes <= VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_bytes;
     -- Outputs
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output := FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output;

     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t[work_inputs_t_bytes_t_h_l69_c45_ff13] LATENCY=0
     -- Inputs
     FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes <= VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes;
     -- Outputs
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output := FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output;

     -- FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t[work_inputs_t_bytes_t_h_l69_c45_ff13] LATENCY=0
     -- Inputs
     FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes <= VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_bytes;
     -- Outputs
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output := FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output;

     -- Submodule level 3
     -- CONST_REF_RD_work_inputs_t_work_inputs_t_1fa3[work_inputs_t_bytes_t_h_l87_c12_d3f7] LATENCY=0
     VAR_CONST_REF_RD_work_inputs_t_work_inputs_t_1fa3_work_inputs_t_bytes_t_h_l87_c12_d3f7_return_output := CONST_REF_RD_work_inputs_t_work_inputs_t_1fa3(
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output,
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_0_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output,
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output,
     VAR_FOR_work_inputs_t_bytes_t_h_l60_c1_7764_ITER_1_FOR_work_inputs_t_bytes_t_h_l62_c1_1d88_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l69_c45_ff13_return_output,
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output,
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_0_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output,
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_0_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output,
     VAR_FOR_work_inputs_t_bytes_t_h_l74_c1_14d0_ITER_1_FOR_work_inputs_t_bytes_t_h_l76_c1_d203_ITER_1_bytes_to_int8_t_work_inputs_t_bytes_t_h_l83_c45_bb36_return_output);

     -- Submodule level 4
     VAR_return_output := VAR_CONST_REF_RD_work_inputs_t_work_inputs_t_1fa3_work_inputs_t_bytes_t_h_l87_c12_d3f7_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
