-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 17
entity work_0CLK_83e31706 is
port(
 inputs : in work_inputs_t;
 return_output : out work_outputs_t);
end work_0CLK_83e31706;
architecture arch of work_0CLK_83e31706 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf]
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS[work_h_l68_c17_2466]
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_right : signed(15 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_return_output : signed(16 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf]
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS[work_h_l68_c17_5cdb]
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_right : signed(15 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_return_output : signed(16 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf]
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS[work_h_l68_c17_daa8]
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_right : signed(15 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_return_output : signed(16 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf]
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS[work_h_l68_c17_8ee7]
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_right : signed(15 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_return_output : signed(16 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf]
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS[work_h_l68_c17_3aa6]
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_right : signed(15 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_return_output : signed(16 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf]
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS[work_h_l68_c17_c097]
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_right : signed(15 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_return_output : signed(16 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf]
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS[work_h_l68_c17_d44c]
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_right : signed(15 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_return_output : signed(16 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf]
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS[work_h_l68_c17_40e2]
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_left : signed(7 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_right : signed(15 downto 0);
signal FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_return_output : signed(16 downto 0);

function CONST_REF_RD_work_outputs_t_work_outputs_t_c871( ref_toks_0 : signed;
 ref_toks_1 : signed;
 ref_toks_2 : signed;
 ref_toks_3 : signed) return work_outputs_t is
 
  variable base : work_outputs_t; 
  variable return_output : work_outputs_t;
begin
      base.result(0)(0) := ref_toks_0;
      base.result(0)(1) := ref_toks_1;
      base.result(1)(0) := ref_toks_2;
      base.result(1)(1) := ref_toks_3;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466 : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_left,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_right,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_left,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_right,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8 : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_left,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_right,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7 : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_left,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_right,
FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6 : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_left,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_right,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097 : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_left,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_right,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_left,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_right,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output);

-- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2 : 0 clocks latency
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_left,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_right,
FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 inputs,
 -- All submodule outputs
 FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output,
 FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_return_output,
 FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output,
 FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_return_output,
 FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output,
 FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_return_output,
 FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output,
 FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_return_output,
 FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output,
 FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_return_output,
 FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output,
 FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_return_output,
 FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output,
 FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_return_output,
 FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output,
 FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : work_outputs_t;
 variable VAR_inputs : work_inputs_t;
 variable VAR_outputs : work_outputs_t;
 variable VAR_i : unsigned(31 downto 0);
 variable VAR_j : unsigned(31 downto 0);
 variable VAR_k : unsigned(31 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_outputs_result_0_0_work_h_l65_c13_d0c8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_0_0_work_h_l68_c17_5711 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_0_0_work_h_l68_c17_5711 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_outputs_result_0_1_work_h_l65_c13_d0c8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_0_1_work_h_l68_c17_5711 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_0_1_work_h_l68_c17_5711 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_outputs_result_1_0_work_h_l65_c13_d0c8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_1_0_work_h_l68_c17_5711 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_1_0_work_h_l68_c17_5711 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_outputs_result_1_1_work_h_l65_c13_d0c8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_1_1_work_h_l68_c17_5711 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_1_1_work_h_l68_c17_5711 : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_return_output : signed(16 downto 0);
 variable VAR_CONST_REF_RD_work_outputs_t_work_outputs_t_c871_work_h_l72_c12_1ca8_return_output : work_outputs_t;
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l68_c41_d2bd_DUPLICATE_03e0_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l68_c64_4b6c_DUPLICATE_040d_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l68_c41_d2bd_DUPLICATE_bce4_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l68_c64_4b6c_DUPLICATE_44a3_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l68_c64_4b6c_DUPLICATE_bb17_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l68_c64_4b6c_DUPLICATE_dbc6_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l68_c41_d2bd_DUPLICATE_21a6_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l68_c41_d2bd_DUPLICATE_c658_return_output : signed(7 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_outputs_result_0_1_work_h_l65_c13_d0c8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_left := VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_outputs_result_0_1_work_h_l65_c13_d0c8;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_outputs_result_1_0_work_h_l65_c13_d0c8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_left := VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_outputs_result_1_0_work_h_l65_c13_d0c8;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_outputs_result_1_1_work_h_l65_c13_d0c8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_left := VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_outputs_result_1_1_work_h_l65_c13_d0c8;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_outputs_result_0_0_work_h_l65_c13_d0c8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_left := VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_outputs_result_0_0_work_h_l65_c13_d0c8;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_inputs := inputs;

     -- Submodule level 0
     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d[work_h_l68_c64_4b6c]_DUPLICATE_040d LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l68_c64_4b6c_DUPLICATE_040d_return_output := VAR_inputs.matrix1(0)(0);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d[work_h_l68_c41_d2bd]_DUPLICATE_bce4 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l68_c41_d2bd_DUPLICATE_bce4_return_output := VAR_inputs.matrix0(0)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d[work_h_l68_c64_4b6c]_DUPLICATE_bb17 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l68_c64_4b6c_DUPLICATE_bb17_return_output := VAR_inputs.matrix1(0)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d[work_h_l68_c41_d2bd]_DUPLICATE_03e0 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l68_c41_d2bd_DUPLICATE_03e0_return_output := VAR_inputs.matrix0(0)(0);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d[work_h_l68_c41_d2bd]_DUPLICATE_c658 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l68_c41_d2bd_DUPLICATE_c658_return_output := VAR_inputs.matrix0(1)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d[work_h_l68_c41_d2bd]_DUPLICATE_21a6 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l68_c41_d2bd_DUPLICATE_21a6_return_output := VAR_inputs.matrix0(1)(0);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d[work_h_l68_c64_4b6c]_DUPLICATE_44a3 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l68_c64_4b6c_DUPLICATE_44a3_return_output := VAR_inputs.matrix1(1)(0);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d[work_h_l68_c64_4b6c]_DUPLICATE_dbc6 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l68_c64_4b6c_DUPLICATE_dbc6_return_output := VAR_inputs.matrix1(1)(1);

     -- Submodule level 1
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l68_c41_d2bd_DUPLICATE_03e0_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l68_c41_d2bd_DUPLICATE_03e0_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l68_c41_d2bd_DUPLICATE_bce4_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l68_c41_d2bd_DUPLICATE_bce4_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l68_c41_d2bd_DUPLICATE_21a6_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l68_c41_d2bd_DUPLICATE_21a6_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l68_c41_d2bd_DUPLICATE_c658_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l68_c41_d2bd_DUPLICATE_c658_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l68_c64_4b6c_DUPLICATE_040d_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l68_c64_4b6c_DUPLICATE_040d_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l68_c64_4b6c_DUPLICATE_bb17_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l68_c64_4b6c_DUPLICATE_bb17_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l68_c64_4b6c_DUPLICATE_44a3_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l68_c64_4b6c_DUPLICATE_44a3_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l68_c64_4b6c_DUPLICATE_dbc6_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l68_c64_4b6c_DUPLICATE_dbc6_return_output;
     -- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left;
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output := FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left;
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output := FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left;
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output := FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left;
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output := FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left;
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output := FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left;
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output := FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left;
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output := FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT[work_h_l68_c41_0caf] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_left;
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output := FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;

     -- Submodule level 2
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_right := VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_right := VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_right := VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_right := VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_right := VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_right := VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_right := VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_right := VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_INFERRED_MULT_work_h_l68_c41_0caf_return_output;
     -- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS[work_h_l68_c17_2466] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_left;
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_return_output := FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS[work_h_l68_c17_daa8] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_left;
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_return_output := FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS[work_h_l68_c17_3aa6] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_left;
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_return_output := FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS[work_h_l68_c17_d44c] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_left;
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_return_output := FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_return_output;

     -- Submodule level 3
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_0_0_work_h_l68_c17_5711 := resize(VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_2466_return_output, 8);
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_0_1_work_h_l68_c17_5711 := resize(VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_daa8_return_output, 8);
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_1_0_work_h_l68_c17_5711 := resize(VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_3aa6_return_output, 8);
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_1_1_work_h_l68_c17_5711 := resize(VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_BIN_OP_PLUS_work_h_l68_c17_d44c_return_output, 8);
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_left := VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_0_0_work_h_l68_c17_5711;
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_left := VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_0_1_work_h_l68_c17_5711;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_left := VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_1_0_work_h_l68_c17_5711;
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_left := VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_0_outputs_result_1_1_work_h_l68_c17_5711;
     -- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS[work_h_l68_c17_c097] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_left;
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_return_output := FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS[work_h_l68_c17_8ee7] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_left;
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_return_output := FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS[work_h_l68_c17_40e2] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_left;
     FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_return_output := FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_return_output;

     -- FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS[work_h_l68_c17_5cdb] LATENCY=0
     -- Inputs
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_left <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_left;
     FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_right <= VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_right;
     -- Outputs
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_return_output := FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_return_output;

     -- Submodule level 4
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_0_0_work_h_l68_c17_5711 := resize(VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_5cdb_return_output, 8);
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_0_1_work_h_l68_c17_5711 := resize(VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_8ee7_return_output, 8);
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_1_0_work_h_l68_c17_5711 := resize(VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_c097_return_output, 8);
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_1_1_work_h_l68_c17_5711 := resize(VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_BIN_OP_PLUS_work_h_l68_c17_40e2_return_output, 8);
     -- CONST_REF_RD_work_outputs_t_work_outputs_t_c871[work_h_l72_c12_1ca8] LATENCY=0
     VAR_CONST_REF_RD_work_outputs_t_work_outputs_t_c871_work_h_l72_c12_1ca8_return_output := CONST_REF_RD_work_outputs_t_work_outputs_t_c871(
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_0_0_work_h_l68_c17_5711,
     VAR_FOR_work_h_l61_c5_fba5_ITER_0_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_0_1_work_h_l68_c17_5711,
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_0_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_1_0_work_h_l68_c17_5711,
     VAR_FOR_work_h_l61_c5_fba5_ITER_1_FOR_work_h_l63_c9_d7e5_ITER_1_FOR_work_h_l66_c13_5760_ITER_1_outputs_result_1_1_work_h_l68_c17_5711);

     -- Submodule level 5
     VAR_return_output := VAR_CONST_REF_RD_work_outputs_t_work_outputs_t_c871_work_h_l72_c12_1ca8_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
